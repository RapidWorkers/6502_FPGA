/*
6502 Implemention in Verilog

Copyright (c) <2019> S.H Kim (soohyunkim@kw.ac.kr)

See the file LICENSE for copying permission.
*/

module BCD_CLA(
    input [7:0] A,//Input A
    input [7:0] B,//Input B
    input Cin,//Carry In
	 output [7:0] S,//BCD Sum
    output Cout,//BCD Carry out
    output HCout//Half Carry Out
);

endmodule
